library verilog;
use verilog.vl_types.all;
entity elevador_rtl_vlg_vec_tst is
end elevador_rtl_vlg_vec_tst;
